`timescale 10 ns/10 ps

module tb();
  
    reg [63:0] in1, in2;
	 reg clk;
	 wire [63:0] out1;
	 
	 reg [63:0] in_data1[0:10];
	 reg [63:0] in_data2[0:10];
	 
	 integer i;
	 
	 initial 
	 begin
	 
	 i = 0;
	 
    in_data1[0] = 64'h4034666666666666;  //-3.14
	 in_data2[0] = 64'hC05891CAC083126F;  //9.2749
	 
	 in_data1[1] = 64'b0100000001001001001001001011110001101010011111101111100111011011;  //50.287
	 in_data2[1] = 64'b0100000001011110000110001011111110110001010110110101011100111111;  //120.3867
	 
	 in_data1[2] = 64'b1100000001011000110010110110111000101110101100011100010000110011;  //-99.1786
	 in_data2[2] = 64'b1100000000000111001011010111011100110001100011111100010100000101;  //-2.8972
	
	 in_data1[3] = 64'b0011111101100101000011011010111000111110011011000100110001011001;  //0.00257
	 in_data2[3] = 64'b0011111111001101010011111101111100111011011001000101101000011101;  //0.229
	 
	 in_data1[4] = 64'b1011111111111110000100000110001001001101110100101111000110101010;  //-1.879
	 in_data2[4] = 64'b1100000000011100111100101011000000100000110001001001101110100110;  //-7.237
	 
	 in_data1[5] = 64'b1011111111101100111010111100010000001000110110001110110010010110;  //-0.90378
	 in_data2[5] = 64'b1100000000011100111100101011000000100000110001001001101110100110;  //-7.237
	 
	 in_data1[6] = 64'b0100000100001000110101101011000111101010011011110011111101010011;  //203478.23947
	 in_data2[6] = 64'b0100000011011000011000111001100101111000110101001111110111110100;  //24974.398
	 
	 in_data1[7] = 64'b1100000001110010000101001010000110101011010010110111001011000101;  //-289.28947
	 in_data2[7] = 64'b1100000010001110011100110010111100011010100111111011111001110111;  //-974.398
	 
	 in_data1[8] = 64'b0100000000101001100100000110001001001101110100101111000110101010;  //12.782
	 in_data2[8] = 64'b0100000001010010011110110101001111110111110011101101100100010111;  //73.927
	 
	 in_data1[9] = 64'b0100000000011001100010010011011101001011110001101010011111110000;  //6.384
	 in_data2[9] = 64'b1100000001011000100100011100101011000000100000110001001001101111;  //-98.278
	 
	 in_data1[10] = 64'b0100000011001000000010000000000000000000000000000000000000000000;  //1234
	 in_data2[10] = 64'b0011111111110000000000000000000000000000000000000000000000000000;  //1
	 
     

	 end

    floating_point_adder UUT (.f_in1(in1), .f_in2(in2), .f_out(out1), .clk(clk));
	 
	 always 
    begin
    clk = 1'b1; 
    #1; // high for 20 * timescale = 20 ns

    clk = 1'b0;
    #1; // low for 20 * timescale = 20 ns
    end 
	
	 always @ (posedge clk)
	 begin
  
	 
	  in1 <= in_data1[i];
	  in2 <= in_data2[i];
	  
	  i = i + 1;
	
    end	
		 
endmodule